magic
tech scmos
magscale 1 3
timestamp 1721563131
<< checkpaint >>
rect -72 -109 96 70
rect -51 -110 96 -109
rect -51 -112 75 -110
<< nwell >>
rect -30 -6 54 69
<< ntransistor >>
rect 9 -69 15 -49
<< ptransistor >>
rect 9 10 15 30
<< ndiffusion >>
rect 6 -69 9 -49
rect 15 -69 18 -49
<< pdiffusion >>
rect 6 10 9 30
rect 15 10 18 30
<< ndcontact >>
rect -12 -69 6 -49
rect 18 -69 36 -49
<< pdcontact >>
rect -12 10 6 30
rect 18 10 36 30
<< psubstratepcontact >>
rect 15 -99 33 -81
<< nsubstratencontact >>
rect 15 42 33 60
<< polysilicon >>
rect 9 30 15 36
rect 9 -49 15 10
rect 9 -75 15 -69
<< polycontact >>
rect -9 -30 9 -9
<< metal1 >>
rect -15 60 36 63
rect -15 42 15 60
rect 33 42 36 60
rect -15 39 36 42
rect -12 30 6 39
rect -15 -30 -9 -9
rect 18 -49 36 10
rect -12 -78 6 -69
rect -15 -81 36 -78
rect -15 -99 15 -81
rect 33 -99 36 -81
rect -15 -102 36 -99
<< labels >>
rlabel metal1 -15 39 15 63 0 vdd
port 2 nsew
rlabel metal1 -15 -102 15 -78 0 gnd
port 3 nsew
rlabel metal1 -15 -30 -9 -9 7 A
port 0 w
rlabel metal1 18 -48 36 9 3 Y
port 1 e
<< end >>