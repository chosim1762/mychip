magic
tech scmos
magscale 1 2
timestamp 1759648187
<< nwell >>
rect -26 1 58 85
<< pwell >>
rect -26 -77 58 1
<< ntransistor >>
rect 13 -29 19 -17
<< ptransistor >>
rect 13 13 19 37
<< ndiffusion >>
rect 10 -29 13 -17
rect 19 -29 22 -17
<< pdiffusion >>
rect 10 13 13 37
rect 19 13 22 37
<< ndcontact >>
rect -2 -29 10 -17
rect 22 -29 34 -17
<< pdcontact >>
rect -2 13 10 37
rect 22 13 34 37
<< psubstratepcontact >>
rect 22 -59 34 -47
<< nsubstratencontact >>
rect 22 55 34 67
<< polysilicon >>
rect 13 37 19 46
rect 13 -17 19 13
rect 13 -38 19 -29
<< polycontact >>
rect 1 -11 13 1
<< metal1 >>
rect -14 67 46 73
rect -14 55 22 67
rect 34 55 46 67
rect -14 49 46 55
rect -2 37 10 49
rect -14 -11 1 1
rect 22 -17 34 13
rect -2 -41 10 -29
rect -14 -47 46 -41
rect -14 -59 22 -47
rect 34 -59 46 -47
rect -14 -65 46 -59
<< labels >>
rlabel metal1 -14 49 46 73 0 vdd
port 28 nsew power bidirectional
rlabel metal1 -14 -65 46 -41 0 gnd
port 14 nsew ground bidirectional
rlabel metal1 -14 -11 1 1 0 Vin
port 1 nsew signal input
<< end >>
