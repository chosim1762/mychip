magic
tech scmos
magscale 1 30
timestamp 1760885258
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal2 >>
rect 43900 48800 46500 49500
<< metal3 >>
rect 80100 145100 80600 146000
rect 92700 145000 93200 146000
rect 107100 144800 107600 146000
rect 121100 144900 121600 146100
rect 144000 139950 145950 140640
rect 144660 122430 146010 123150
rect 144660 109740 145950 110040
rect 144800 94200 145900 94600
rect 144500 64400 146000 64800
rect 144700 58700 146200 59100
rect 50300 44000 50800 45400
rect 64700 44100 65200 45300
rect 90000 43800 90700 45800
rect 115900 44100 116400 44900
rect 130900 44100 131500 44500
<< end >>