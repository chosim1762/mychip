magic
tech scmos
timestamp 1759672588
<< nwell >>
rect -16 3 14 34
<< pwell >>
rect -16 -33 14 3
<< ntransistor >>
rect -2 -20 0 -14
<< ptransistor >>
rect -2 9 0 21
<< ndiffusion >>
rect -4 -20 -2 -14
rect 0 -20 2 -14
<< pdiffusion >>
rect -4 9 -2 21
rect 0 9 2 21
<< ndcontact >>
rect -10 -20 -4 -14
rect 2 -20 8 -14
<< pdcontact >>
rect -10 9 -4 21
rect 2 9 8 21
<< psubstratepcontact >>
rect 1 -30 7 -24
<< nsubstratencontact >>
rect 2 25 8 31
<< polysilicon >>
rect -2 21 0 23
rect -2 1 0 9
rect -2 -14 0 -5
rect -2 -22 0 -20
<< polycontact >>
rect -7 -5 0 1
<< metal1 >>
rect -13 25 2 31
rect 8 25 11 31
rect -10 21 -4 25
rect -11 -5 -7 1
rect 8 -20 11 21
rect -10 -24 -4 -20
rect -11 -30 1 -24
rect 7 -30 10 -24
<< labels >>
rlabel metal1 -13 25 2 31 0 vdd
port 1 nsew
rlabel metal1 -11 -30 1 -24 0 gnd
port 2 nsew
rlabel metal1 -11 -5 0 1 0 Vin
port 1 nsew signal input
rlabel metal1 8 -20 11 21 0 Vout
port 2 nsew signal output
<< end >>
