magic
tech scmos
magscale 1 4
timestamp 1760883564
<< checkpaint >>
rect 10680 19290 10880 19544
rect 12360 19264 12560 19544
rect 14280 19238 14480 19544
rect 16144 19251 16344 19544
rect 19238 18560 19544 18784
rect 19316 16224 19544 16440
rect 19290 14520 19544 14720
rect 19316 12452 19544 12652
rect 19277 8480 19544 8680
rect 19290 7720 19544 7920
rect 5784 6412 6294 6640
rect 6704 5784 6904 6073
rect 8624 5784 8824 6047
rect 12012 5784 12224 6099
rect 15440 5784 15640 6008
<< nwell >>
rect 16680 8980 16828 9136
rect 18292 8940 18544 9096
rect 6920 7336 7196 7540
rect 15824 7324 16072 7500
rect 8864 7144 8984 7268
rect 12264 7104 12400 7228
rect 17668 7168 18004 7504
<< pwell >>
rect 18292 8800 18544 8940
rect 6920 6904 7196 7336
rect 8864 7000 8984 7144
rect 12264 6960 12400 7104
rect 15824 7012 16072 7324
rect 17668 6856 18004 7168
<< ntransistor >>
rect 16760 8872 16772 8904
rect 18408 8860 18416 8884
rect 15912 7152 15932 7188
rect 7008 7056 7040 7100
rect 8920 7052 8928 7076
rect 17824 7048 17848 7096
rect 12328 7012 12336 7036
<< ptransistor >>
rect 16760 9020 16772 9036
rect 18408 8968 18416 9012
rect 7016 7376 7036 7408
rect 15912 7372 15932 7404
rect 8920 7168 8928 7216
rect 17824 7216 17848 7312
rect 12328 7128 12336 7176
<< ndiffusion >>
rect 16752 8872 16760 8904
rect 16772 8872 16780 8904
rect 18404 8860 18408 8884
rect 18416 8860 18420 8884
rect 15908 7152 15912 7188
rect 15932 7152 15936 7188
rect 7000 7056 7008 7100
rect 7040 7056 7048 7100
rect 7088 7056 7092 7100
rect 8912 7052 8920 7076
rect 8928 7052 8936 7076
rect 17812 7048 17824 7096
rect 17848 7048 17860 7096
rect 12316 7012 12328 7036
rect 12336 7012 12348 7036
<< pdiffusion >>
rect 16752 9020 16760 9036
rect 16772 9020 16780 9036
rect 18392 8968 18408 9012
rect 18416 8968 18432 9012
rect 7004 7376 7016 7408
rect 7036 7376 7048 7408
rect 15908 7372 15912 7404
rect 15932 7372 15936 7404
rect 8912 7168 8920 7216
rect 8928 7168 8936 7216
rect 17812 7216 17824 7312
rect 17848 7216 17860 7312
rect 12316 7128 12328 7176
rect 12336 7128 12348 7176
<< ndcontact >>
rect 16728 8872 16752 8904
rect 16780 8872 16804 8904
rect 18364 8860 18404 8884
rect 18420 8860 18460 8884
rect 15876 7152 15908 7188
rect 15936 7152 15968 7188
rect 6960 7056 7000 7100
rect 7048 7056 7088 7100
rect 8888 7052 8912 7076
rect 8936 7052 8960 7076
rect 15964 7048 15996 7080
rect 17764 7048 17812 7096
rect 17860 7048 17908 7096
rect 12288 7012 12316 7036
rect 12348 7012 12376 7036
rect 7084 6936 7116 6968
<< pdcontact >>
rect 16728 9008 16752 9036
rect 16780 9008 16804 9036
rect 18364 8968 18392 9012
rect 18432 8968 18460 9012
rect 7096 7476 7128 7508
rect 6972 7376 7004 7408
rect 7048 7376 7080 7408
rect 15876 7372 15908 7404
rect 15936 7372 15968 7404
rect 8888 7168 8912 7216
rect 8936 7168 8960 7216
rect 17764 7216 17812 7312
rect 17860 7216 17908 7312
rect 12288 7128 12316 7176
rect 12348 7128 12376 7176
<< psubstratepcontact >>
rect 16768 8816 16792 8840
rect 18412 8812 18436 8836
rect 8932 7012 8956 7036
rect 12348 6968 12372 6996
rect 17860 6928 17908 6976
<< nsubstratencontact >>
rect 16768 9056 16796 9088
rect 18408 9032 18432 9056
rect 17860 7384 17908 7432
rect 8936 7232 8960 7256
rect 12352 7192 12376 7220
<< polysilicon >>
rect 16760 9036 16772 9044
rect 16760 8904 16772 9020
rect 18408 9012 18416 9020
rect 18408 8928 18416 8968
rect 18408 8884 18416 8904
rect 16760 8860 16772 8872
rect 18408 8852 18416 8860
rect 7016 7408 7036 7432
rect 15912 7404 15932 7420
rect 7016 7364 7036 7376
rect 15912 7348 15932 7372
rect 17824 7312 17848 7348
rect 8920 7216 8928 7224
rect 15912 7188 15932 7220
rect 12328 7176 12336 7184
rect 8920 7136 8928 7168
rect 7008 7100 7040 7116
rect 15912 7136 15932 7152
rect 8920 7076 8928 7112
rect 12328 7112 12336 7128
rect 12328 7096 12336 7104
rect 17824 7096 17848 7216
rect 7008 7044 7040 7056
rect 8920 7044 8928 7052
rect 12328 7036 12336 7072
rect 17824 7012 17848 7048
rect 12328 7004 12336 7012
<< polycontact >>
rect 16736 8928 16760 8956
rect 18400 8904 18424 8928
rect 7000 7316 7052 7364
rect 15904 7312 15940 7348
rect 15904 7220 15940 7256
rect 6996 7116 7052 7168
rect 8900 7112 8928 7136
rect 17776 7120 17824 7168
rect 12328 7104 12336 7112
<< metal1 >>
rect 10744 19240 10812 19252
rect 10744 19200 10760 19240
rect 10800 19200 10812 19240
rect 10744 16984 10812 19200
rect 12424 19200 12492 19212
rect 12424 19160 12440 19200
rect 12480 19160 12492 19200
rect 12424 17492 12492 19160
rect 14344 19160 14412 19172
rect 14344 19120 14360 19160
rect 14400 19120 14412 19160
rect 14344 19104 14412 19120
rect 16200 19160 16292 19184
rect 16200 19104 16224 19160
rect 16264 19104 16292 19160
rect 14360 17892 14400 19104
rect 14344 17880 14412 17892
rect 14344 17840 14360 17880
rect 14400 17840 14412 17880
rect 14344 17824 14412 17840
rect 12424 17452 12440 17492
rect 12480 17452 12492 17492
rect 12424 17440 12492 17452
rect 10744 16944 10760 16984
rect 10800 16944 10812 16984
rect 10744 16932 10812 16944
rect 12572 16344 12640 16360
rect 12572 16304 12584 16344
rect 12624 16304 12640 16344
rect 12572 16292 12640 16304
rect 9092 14640 9160 14652
rect 9092 14600 9104 14640
rect 9144 14600 9160 14640
rect 9092 14584 9160 14600
rect 7344 12572 7440 12600
rect 7344 12532 7372 12572
rect 7412 12532 7440 12572
rect 7344 12504 7440 12532
rect 7080 7960 7144 8024
rect 7092 7532 7132 7960
rect 7080 7512 7144 7532
rect 6956 7508 7176 7512
rect 6956 7476 7096 7508
rect 7128 7476 7176 7508
rect 6956 7472 7176 7476
rect 6968 7408 7004 7472
rect 7080 7464 7144 7472
rect 6968 7376 6972 7408
rect 7080 7376 7168 7408
rect 7000 7312 7052 7316
rect 6996 7264 7052 7312
rect 6772 7216 7052 7264
rect 7124 7252 7168 7376
rect 7372 7252 7412 12504
rect 8880 7904 8944 7920
rect 8880 7864 8892 7904
rect 8932 7864 8944 7904
rect 8880 7852 8944 7864
rect 8892 7256 8932 7852
rect 6772 7212 6960 7216
rect 6772 7052 6840 7212
rect 6996 7168 7052 7216
rect 7120 7212 7412 7252
rect 8876 7232 8936 7256
rect 8960 7232 8972 7256
rect 8888 7216 8912 7232
rect 6772 6132 6784 7052
rect 6824 6132 6840 7052
rect 6956 7100 7000 7104
rect 7124 7100 7168 7212
rect 8960 7144 8972 7216
rect 9104 7144 9144 14584
rect 12292 7944 12360 7960
rect 12292 7904 12304 7944
rect 12344 7904 12360 7944
rect 12292 7892 12360 7904
rect 12304 7220 12344 7892
rect 12276 7192 12352 7220
rect 12376 7192 12388 7220
rect 6956 7056 6960 7100
rect 7000 7056 7048 7100
rect 7088 7056 7168 7100
rect 8692 7136 8892 7144
rect 8692 7112 8900 7136
rect 8692 7104 8892 7112
rect 8960 7104 9144 7144
rect 12288 7176 12316 7192
rect 12092 7112 12320 7120
rect 12092 7104 12328 7112
rect 12376 7104 12388 7176
rect 12584 7104 12624 16292
rect 15944 7904 16012 7920
rect 15944 7864 15960 7904
rect 16000 7864 16012 7904
rect 15944 7852 16012 7864
rect 15960 7468 16000 7852
rect 15860 7440 16036 7468
rect 15876 7404 15908 7440
rect 15904 7304 15940 7312
rect 6956 6972 7000 7056
rect 7064 6972 7132 6984
rect 6956 6968 7132 6972
rect 6956 6936 7084 6968
rect 7116 6936 7132 6968
rect 6956 6932 7132 6936
rect 7064 6920 7132 6932
rect 7080 6852 7120 6920
rect 7064 6840 7132 6852
rect 7064 6800 7080 6840
rect 7120 6800 7132 6840
rect 7064 6784 7132 6800
rect 6772 6120 6840 6132
rect 6772 6080 6784 6120
rect 6824 6080 6840 6120
rect 8692 6144 8760 7104
rect 8960 7052 8972 7104
rect 12092 7092 12320 7104
rect 8888 7036 8912 7052
rect 8884 7012 8932 7036
rect 8956 7012 8968 7036
rect 8892 6944 8932 7012
rect 8880 6932 8944 6944
rect 8880 6892 8892 6932
rect 8932 6892 8944 6932
rect 8880 6880 8944 6892
rect 12092 6240 12144 7092
rect 12376 7064 12624 7104
rect 15520 7264 15940 7304
rect 12376 7012 12388 7064
rect 12288 6996 12316 7012
rect 12284 6968 12348 6996
rect 12372 6968 12384 6996
rect 12304 6892 12344 6968
rect 12292 6880 12360 6892
rect 12292 6840 12304 6880
rect 12344 6840 12360 6880
rect 12292 6824 12360 6840
rect 12080 6224 12160 6240
rect 12080 6172 12092 6224
rect 12144 6172 12160 6224
rect 12080 6160 12160 6172
rect 8692 6104 8704 6144
rect 8744 6104 8760 6144
rect 8692 6092 8760 6104
rect 6772 6064 6840 6080
rect 15520 6052 15560 7264
rect 15904 7256 15940 7264
rect 15968 7320 16000 7408
rect 16200 7320 16212 19104
rect 15968 7304 16212 7320
rect 15968 7240 15984 7304
rect 16280 7240 16292 19104
rect 17984 17880 18052 17892
rect 17984 17840 18000 17880
rect 18040 17840 18052 17880
rect 17012 17492 17080 17504
rect 17012 17452 17024 17492
rect 17064 17452 17080 17492
rect 17012 17440 17080 17452
rect 16704 9224 16772 9240
rect 16704 9184 16720 9224
rect 16760 9184 16772 9224
rect 16704 9172 16772 9184
rect 16720 9092 16760 9172
rect 16720 9088 16816 9092
rect 16720 9080 16768 9088
rect 16724 9056 16768 9080
rect 16796 9056 16816 9088
rect 16724 9052 16816 9056
rect 16728 9036 16752 9052
rect 16780 8960 16804 9008
rect 17024 8960 17064 17440
rect 16504 8956 16732 8960
rect 16504 8928 16736 8956
rect 16504 8920 16732 8928
rect 16780 8920 17064 8960
rect 16504 7852 16572 8920
rect 16780 8904 16804 8920
rect 16728 8844 16752 8872
rect 16724 8840 16816 8844
rect 16724 8824 16768 8840
rect 16720 8816 16768 8824
rect 16792 8816 16816 8840
rect 16720 8812 16816 8816
rect 16720 8664 16760 8812
rect 16692 8640 16784 8664
rect 16692 8600 16720 8640
rect 16760 8600 16784 8640
rect 16692 8572 16784 8600
rect 17744 8040 17812 8052
rect 17744 8000 17760 8040
rect 17800 8000 17812 8040
rect 17744 7984 17812 8000
rect 16504 7812 16520 7852
rect 16560 7812 16572 7852
rect 16504 7800 16572 7812
rect 17760 7456 17800 7984
rect 17716 7432 17956 7456
rect 17716 7384 17860 7432
rect 17908 7384 17956 7432
rect 17716 7360 17956 7384
rect 17760 7312 17812 7360
rect 17760 7292 17764 7312
rect 15968 7224 16292 7240
rect 15968 7152 16000 7224
rect 17860 7184 17908 7216
rect 17984 7184 18052 17840
rect 18172 16984 18240 17000
rect 18172 16944 18184 16984
rect 18224 16944 18240 16984
rect 18172 16932 18240 16944
rect 18184 9600 18224 16932
rect 18492 16344 18560 16360
rect 19240 16344 19304 16360
rect 18492 16304 18504 16344
rect 18544 16304 19252 16344
rect 19292 16304 19304 16344
rect 18492 16292 18560 16304
rect 19240 16292 19304 16304
rect 18480 14640 19292 14652
rect 18480 14600 18492 14640
rect 18532 14600 19240 14640
rect 19280 14600 19292 14640
rect 18480 14584 19292 14600
rect 18532 12584 18624 12600
rect 18532 12520 18544 12584
rect 18612 12572 18624 12584
rect 19224 12572 19320 12600
rect 18612 12532 19252 12572
rect 19292 12532 19320 12572
rect 18612 12520 18624 12532
rect 18532 12504 18624 12520
rect 19224 12504 19320 12532
rect 18184 9560 18664 9600
rect 18332 9240 18424 9252
rect 18332 9172 18344 9240
rect 18412 9172 18424 9240
rect 18332 9160 18424 9172
rect 18360 9060 18400 9160
rect 18356 9056 18436 9060
rect 18356 9032 18408 9056
rect 18432 9032 18436 9056
rect 18356 9028 18436 9032
rect 18364 9012 18392 9028
rect 18460 8932 18472 9012
rect 18624 8932 18664 9560
rect 18160 8928 18384 8932
rect 18160 8904 18400 8928
rect 18160 8892 18384 8904
rect 18460 8892 18664 8932
rect 18160 8612 18212 8892
rect 18460 8860 18472 8892
rect 18364 8844 18404 8860
rect 18364 8836 18440 8844
rect 18364 8812 18412 8836
rect 18436 8812 18440 8836
rect 18160 8572 18172 8612
rect 18160 8560 18212 8572
rect 18360 8804 18440 8812
rect 18360 8464 18400 8804
rect 18520 8600 18584 8612
rect 19212 8600 19280 8612
rect 18520 8560 18532 8600
rect 18572 8560 19224 8600
rect 19264 8560 19280 8600
rect 18520 8544 18584 8560
rect 19212 8544 19280 8560
rect 18344 8452 18412 8464
rect 18344 8412 18360 8452
rect 18400 8412 18412 8452
rect 18344 8400 18412 8412
rect 18332 7840 18400 7852
rect 19212 7840 19280 7852
rect 18332 7800 18344 7840
rect 18384 7800 19224 7840
rect 19264 7800 19280 7840
rect 18332 7784 18400 7800
rect 19212 7784 19280 7800
rect 17532 7168 17760 7172
rect 17812 7168 18052 7184
rect 15876 7084 15908 7152
rect 17532 7132 17776 7168
rect 15860 7080 16020 7084
rect 15860 7048 15964 7080
rect 15996 7048 16020 7080
rect 15860 7044 16020 7048
rect 15904 6920 15944 7044
rect 15892 6904 15960 6920
rect 15892 6864 15904 6904
rect 15944 6864 15960 6904
rect 15892 6852 15960 6864
rect 15504 6040 15572 6052
rect 15504 6000 15520 6040
rect 15560 6000 15572 6040
rect 17532 6012 17572 7132
rect 17716 7120 17776 7132
rect 17824 7144 18052 7168
rect 17860 7096 17908 7144
rect 17760 7048 17764 7052
rect 17760 7000 17812 7048
rect 17716 6976 17956 7000
rect 17716 6928 17860 6976
rect 17908 6928 17956 6976
rect 17716 6904 17956 6928
rect 17760 6892 17800 6904
rect 17744 6880 17812 6892
rect 17744 6840 17760 6880
rect 17800 6840 17812 6880
rect 17744 6824 17812 6840
rect 15504 5984 15572 6000
rect 17520 6000 17584 6012
rect 17520 5960 17532 6000
rect 17572 5960 17584 6000
rect 17520 5944 17584 5960
<< rmetal1 >>
rect 16224 19104 16264 19120
rect 6784 6132 6824 7052
rect 16212 7304 16280 19104
rect 15984 7240 16280 7304
rect 18544 12572 18612 12584
rect 18544 12532 18560 12572
rect 18600 12532 18612 12572
rect 18544 12520 18612 12532
rect 18344 9224 18412 9240
rect 18344 9184 18360 9224
rect 18400 9184 18412 9224
rect 18344 9172 18412 9184
<< m2contact >>
rect 10760 19200 10800 19240
rect 12440 19160 12480 19200
rect 14360 19120 14400 19160
rect 16224 19120 16264 19160
rect 14360 17840 14400 17880
rect 12440 17452 12480 17492
rect 10760 16944 10800 16984
rect 12584 16304 12624 16344
rect 9104 14600 9144 14640
rect 7372 12532 7412 12572
rect 8892 7864 8932 7904
rect 12304 7904 12344 7944
rect 15960 7864 16000 7904
rect 7080 6800 7120 6840
rect 6784 6080 6824 6120
rect 8892 6892 8932 6932
rect 12304 6840 12344 6880
rect 12092 6172 12144 6224
rect 8704 6104 8744 6144
rect 18000 17840 18040 17880
rect 17024 17452 17064 17492
rect 16720 9184 16760 9224
rect 16720 8600 16760 8640
rect 17760 8000 17800 8040
rect 16520 7812 16560 7852
rect 18184 16944 18224 16984
rect 18504 16304 18544 16344
rect 19252 16304 19292 16344
rect 18492 14600 18532 14640
rect 19240 14600 19280 14640
rect 18560 12532 18600 12572
rect 19252 12532 19292 12572
rect 18360 9184 18400 9224
rect 18172 8572 18212 8612
rect 18532 8560 18572 8600
rect 19224 8560 19264 8600
rect 18360 8412 18400 8452
rect 18344 7800 18384 7840
rect 19224 7800 19264 7840
rect 15904 6864 15944 6904
rect 15520 6000 15560 6040
rect 17760 6840 17800 6880
rect 17532 5960 17572 6000
<< metal2 >>
rect 6464 18840 6532 18852
rect 6464 18800 6480 18840
rect 6520 18800 6532 18840
rect 6464 9384 6532 18800
rect 18864 18840 18932 18852
rect 18864 18800 18880 18840
rect 18920 18800 18932 18840
rect 6612 18692 18784 18704
rect 6612 18652 6624 18692
rect 6664 18652 18732 18692
rect 18772 18652 18784 18692
rect 6612 18640 18784 18652
rect 9092 14640 9160 14652
rect 9092 14600 9104 14640
rect 9144 14600 9160 14640
rect 9092 14584 9160 14600
rect 18864 9384 18932 18800
rect 6464 9320 18932 9384
rect 6464 8172 6532 9320
rect 16720 9252 16760 9320
rect 18360 9252 18400 9320
rect 16692 9224 16784 9252
rect 16692 9184 16720 9224
rect 16760 9184 16784 9224
rect 16692 9160 16784 9184
rect 18332 9224 18424 9252
rect 18332 9184 18360 9224
rect 18400 9184 18424 9224
rect 18332 9160 18424 9184
rect 18864 8172 18932 9320
rect 6464 8104 18932 8172
rect 6464 6560 6532 8104
rect 7092 8024 7132 8104
rect 7080 8012 7144 8024
rect 7080 7972 7092 8012
rect 7132 7972 7144 8012
rect 7080 7960 7144 7972
rect 8892 7920 8932 8104
rect 12304 7960 12344 8104
rect 12292 7944 12360 7960
rect 8880 7904 8944 7920
rect 8880 7864 8892 7904
rect 8932 7864 8944 7904
rect 12292 7904 12304 7944
rect 12344 7904 12360 7944
rect 15960 7932 16000 8104
rect 17760 8052 17800 8104
rect 17744 8040 17812 8052
rect 17744 8000 17760 8040
rect 17800 8000 17812 8040
rect 17744 7984 17812 8000
rect 12292 7892 12360 7904
rect 15932 7904 16024 7932
rect 8880 7852 8944 7864
rect 15932 7864 15960 7904
rect 16000 7864 16024 7904
rect 15932 7840 16024 7864
rect 8880 6932 8944 6944
rect 8880 6892 8892 6932
rect 8932 6892 8944 6932
rect 15880 6904 15972 6932
rect 8880 6880 8944 6892
rect 12292 6880 12360 6892
rect 7064 6840 7132 6852
rect 7064 6800 7080 6840
rect 7120 6800 7132 6840
rect 7064 6784 7132 6800
rect 7080 6704 7120 6784
rect 8892 6704 8932 6880
rect 12292 6840 12304 6880
rect 12344 6840 12360 6880
rect 15880 6864 15904 6904
rect 15944 6864 15972 6904
rect 15880 6840 15972 6864
rect 17744 6880 17812 6892
rect 17744 6840 17760 6880
rect 17800 6840 17812 6880
rect 12292 6824 12360 6840
rect 12304 6704 12344 6824
rect 15904 6704 15944 6840
rect 17744 6824 17812 6840
rect 17760 6704 17800 6824
rect 6612 6692 18784 6704
rect 6612 6652 6624 6692
rect 6664 6652 18732 6692
rect 18772 6652 18784 6692
rect 6612 6640 18784 6652
rect 6214 6544 6532 6560
rect 6214 6504 6480 6544
rect 6520 6504 6532 6544
rect 6214 6492 6532 6504
rect 18864 6544 18932 8104
rect 18864 6504 18880 6544
rect 18920 6504 18932 6544
rect 18864 6492 18932 6504
<< m3contact >>
rect 6480 18800 6520 18840
rect 18880 18800 18920 18840
rect 6624 18652 6664 18692
rect 18732 18652 18772 18692
rect 7092 7972 7132 8012
rect 6624 6652 6664 6692
rect 18732 6652 18772 6692
rect 6480 6504 6520 6544
rect 18880 6504 18920 6544
<< metal3 >>
rect 10760 19264 10800 19370
rect 10732 19184 10824 19264
rect 12440 19212 12480 19344
rect 12424 19144 12492 19212
rect 14360 19172 14400 19318
rect 16224 19184 16264 19331
rect 14344 19104 14412 19172
rect 16200 19092 16292 19184
rect 6464 18840 18932 18852
rect 6464 18800 6480 18840
rect 6520 18800 18880 18840
rect 18920 18800 18932 18840
rect 6464 18784 18932 18800
rect 6612 18692 6680 18704
rect 6612 18652 6624 18692
rect 6664 18652 6680 18692
rect 6612 8332 6680 18652
rect 18720 18692 19318 18704
rect 18720 18652 18732 18692
rect 18772 18652 19318 18692
rect 18720 18640 19318 18652
rect 14344 17880 14412 17892
rect 17984 17880 18052 17892
rect 14344 17840 18052 17880
rect 14344 17824 14412 17840
rect 17984 17824 18052 17840
rect 12412 17492 12504 17520
rect 17000 17492 17092 17520
rect 12412 17452 17092 17492
rect 12412 17424 12504 17452
rect 17000 17424 17092 17452
rect 10732 16984 10824 17012
rect 18160 16984 18252 17012
rect 10732 16944 18252 16984
rect 10732 16920 10824 16944
rect 18160 16920 18252 16944
rect 12572 16344 12640 16360
rect 18480 16344 18572 16372
rect 12572 16304 18572 16344
rect 12572 16292 12640 16304
rect 18480 16280 18572 16304
rect 18464 14640 18560 14664
rect 9160 14600 18560 14640
rect 18464 14572 18560 14600
rect 7344 12572 7440 12600
rect 18532 12572 18624 12600
rect 7344 12532 18624 12572
rect 7344 12504 7440 12532
rect 18532 12504 18624 12532
rect 16692 8572 16784 8664
rect 18144 8600 18224 8612
rect 18504 8600 18600 8624
rect 16720 8332 16760 8572
rect 18144 8560 18600 8600
rect 18144 8544 18224 8560
rect 18504 8532 18600 8560
rect 18332 8384 18424 8480
rect 18360 8332 18400 8384
rect 18720 8332 18784 18640
rect 19224 16360 19320 16372
rect 19224 16304 19396 16360
rect 19224 16280 19320 16304
rect 19212 14640 19304 14664
rect 19212 14600 19370 14640
rect 19212 14572 19304 14600
rect 19224 12572 19320 12600
rect 19224 12532 19396 12572
rect 19224 12504 19320 12532
rect 19200 8600 19292 8624
rect 19200 8560 19357 8600
rect 19200 8532 19292 8560
rect 6612 8264 18784 8332
rect 6612 6692 6680 8264
rect 16492 7840 16584 7864
rect 18320 7840 18412 7864
rect 16492 7800 18412 7840
rect 16492 7784 16584 7800
rect 18320 7772 18412 7800
rect 6612 6652 6624 6692
rect 6664 6652 6680 6692
rect 6612 6640 6680 6652
rect 18720 6692 18784 8264
rect 19200 7840 19292 7864
rect 19200 7800 19370 7840
rect 19200 7772 19292 7800
rect 18720 6652 18732 6692
rect 18772 6652 18784 6692
rect 18720 6640 18784 6652
rect 6464 6544 18932 6560
rect 6464 6504 6480 6544
rect 6520 6504 18880 6544
rect 18920 6504 18932 6544
rect 6464 6492 18932 6504
rect 6760 6052 6852 6144
rect 8680 6080 8772 6160
rect 12064 6144 12172 6252
rect 6784 5993 6824 6052
rect 8704 5967 8744 6080
rect 12092 6019 12144 6144
rect 15492 5972 15584 6064
rect 15520 5928 15560 5972
rect 17504 5932 17600 6024
rect 17532 5864 17572 5932
<< labels >>
rlabel space 6786 5993 6825 6045 0 Vi_G
port 1 nsew
rlabel metal2 6240 6500 6422 6552 1 vdd
port 2 n
rlabel metal3 8710 5980 8736 6045 0 Vi_C
port 3 nsew
rlabel metal3 12103 6032 12142 6097 0 Vi_B
port 4 nsew
rlabel space 15522 5928 15561 5967 0 Vi_A
port 5 nsew
rlabel space 17537 5876 17576 5915 0 Vi_F
port 6 nsew
rlabel metal3 19292 7800 19370 7839 0 Vi_D
port 7 nsew
rlabel metal3 19305 8567 19357 8593 0 Vi_E
port 8 nsew
rlabel space 19396 12506 19474 12584 0 Vo_G
port 9 nsew
rlabel space 19305 14599 19357 14638 0 Vo_C
port 10 nsew
rlabel space 19331 16302 19383 16354 0 Vo_B
port 11 nsew
rlabel space 19149 18642 19305 18707 0 gnd
port 12 nsew
rlabel metal3 16224 19214 16263 19318 0 Vo_A
port 13 nsew
rlabel space 14352 19188 14404 19318 0 Vo_F
port 14 nsew
rlabel metal3 12441 19227 12480 19331 0 Vo_D
port 15 nsew
rlabel space 10764 19279 10803 19357 0 Vo_E
port 16 nsew
<< end >>
